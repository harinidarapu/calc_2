// Transaction class
// Creating randam bit to inputs
//
//          		----------------
//  Port A 			|				|
//req_A [0:3]  -->	|               |  -->out_res_A [0:1]
//Data_A1[0:31]-->	|               |  -->out_Data_A [0:31]
//Data_A2[0:31]  	|               |  -->out_tag_A [0:1]
//tag_A[0:1]   --> 	|               |
//					|               |
//					|               |
//					|               |
//					-----------------

// Similarly we have port A, port B, Port C, Port D

class Transaction
// defining all inputs portwise

	rand bit [0:3] req_A,req_B,req_C,req_D;
	rand bit [0:31] data_A1,data_A2,data_B1,data_B2,data_C1,data_C2,data_D1,data_D2;
	//out_Data_A,out_Data_B,out_Data_C,out_Data_D;
	randc bit [0:1] tag_A,tag_B,tag_C,tag_D;
	bit reset;
	
// puting constraint on the randomly generated stimulus
	constraint req {req_A inside {0,1,2,5,6};
					req_B inside {0,1,2,5,6};
					req_C inside {0,1,2,5,6};
					req_D inside {0,1,2,5,6};
					}
//Print the values generated by transaction class

  function void print_transaction(string class_name);
   		$display ($time," : %s PORTA opcode : %d  data_A1 : %h data_A2 : %h	tag: %h",class_name,req_A,data_A1,data_A2,tag_A );
		$display ($time," : %s PORTB opcode : %d  data_B1 : %h data_B2 : %h	tag: %h",class_name,req_B,data_B1,data_B2,tag_B);
		$display ($time," : %s PORTC opcode : %d  data_C1 : %h data_C2 : %h	tag: %h",class_name,req_C,data_C1,data_C2,tag_C );
		$display ($time," : %s PORTD opcode : %d  data_D1 : %h data_D2: %h	tag: %h",class_name,req_D,data_D1,data_D2,tag_D );
	endfunction: print_transaction
	
endclass